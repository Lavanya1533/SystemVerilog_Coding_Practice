// File name   : counter_test.sv
