// Project     : SystemVerilog Training
